module pipe_ex2(Zout,rs1,rs2,rd,func,addr,clk1,clk2);
endmodule
